`timescale 1ns/1ps
`include "../hdl/defines.v"

module tb_my_riscv ();
    reg r_Clk;
    reg r_reset;
    reg r_ce;
    
    parameter CLK_PERIOD = 40;

endmodule
